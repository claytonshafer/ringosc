* ELDO netlist generated with ICnet by 'cms156' on Tue Mar  8 2022 at 16:34:50

.CONNECT GROUND 0

*
* Globals.
*
.global VDD VSS GROUND

*
* Component pathname : $GDKGATES/inv01
*
.subckt INV01  Y A VDD_ESC1 VSS_ESC2

        MP1 Y A VDD_ESC1 VDD_ESC1 pmos w=0.77u l=0.14u m=1 as=0.2618p ad=0.2618p
+  ps=1.45u pd=1.45u
        MN1 Y A VSS_ESC2 VSS_ESC2 nmos w=0.35u l=0.14u m=1 as=0.119p ad=0.119p
+  ps=1.03u pd=1.03u
.ends INV01

*
* MAIN CELL: Component pathname : $PROJ/ringosc/rlc
*
        X_INV014 N$69 N$71 VDD VSS INV01
        X_INV015 N$71 OUT VDD VSS INV01
        X_INV012 N$64 N$70 VDD VSS INV01
        X_INV013 N$70 N$69 VDD VSS INV01
        X_INV011 OUT N$64 VDD VSS INV01
        V1 N$13 GROUND DC 5V
        V2 VSS GROUND DC 0V
        R1 N$13 N$55 200 NOISE=1
        C1 VDD VSS 100p
        L1 N$55 VDD 0.1u
*
.end
